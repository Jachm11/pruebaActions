// Simple AND gate module in Verilog

module and_gate 

(
          input  wire a,  // First input
input  wire b  // Second input 
);
      assign y = a & b;  // Output is the AND of inputs a and b










    endmodule